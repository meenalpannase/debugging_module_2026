// =========================================================================
  // SPI AGENT
  // =========================================================================
  
  class spi_agent extends uvm_agent;
    `uvm_component_utils(spi_agent)
    
    spi_driver    driver;
    spi_monitor   monitor;
    spi_sequencer sequencer;
    spi_config    cfg;
    
    uvm_analysis_port #(spi_transaction) analysis_port;
    
    function new(string name, uvm_component parent);
      super.new(name, parent);
    endfunction
    
    virtual function void build_phase(uvm_phase phase);
      super.build_phase(phase);
      
      if (!uvm_config_db#(spi_config)::get(this, "", "cfg", cfg))
        `uvm_fatal(get_type_name(), "Config not found")
      
      monitor = spi_monitor::type_id::create("monitor", this);
      
      if (cfg.is_active == UVM_ACTIVE) begin
        driver = spi_driver::type_id::create("driver", this);
        sequencer = spi_sequencer::type_id::create("sequencer", this);
      end
    endfunction
    
    virtual function void connect_phase(uvm_phase phase);
      super.connect_phase(phase);
      
      if (cfg.is_active == UVM_ACTIVE) begin
        driver.seq_item_port.connect(sequencer.seq_item_export);
      end
      
      analysis_port = monitor.analysis_port;
    endfunction
    
  endclass
  
